module halfadder (input a, b,
                  output s, c);

endmodule // halfadder
